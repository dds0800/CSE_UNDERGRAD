library verilog;
use verilog.vl_types.all;
entity Overflow_vlg_check_tst is
    port(
        OVER            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Overflow_vlg_check_tst;
