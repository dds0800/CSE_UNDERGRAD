library verilog;
use verilog.vl_types.all;
entity ALUXOR_vlg_vec_tst is
end ALUXOR_vlg_vec_tst;
