library verilog;
use verilog.vl_types.all;
entity Overflow_vlg_vec_tst is
end Overflow_vlg_vec_tst;
