library verilog;
use verilog.vl_types.all;
entity AdderSubtractor_vlg_vec_tst is
end AdderSubtractor_vlg_vec_tst;
