library verilog;
use verilog.vl_types.all;
entity ALUAND_vlg_vec_tst is
end ALUAND_vlg_vec_tst;
